--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   03:10:34 03/23/2025
-- Design Name:   
-- Module Name:   /home/ise/vhdl/DeMuX_1_4/DeMuX_1_4_TB.vhd
-- Project Name:  DeMuX_1_4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: DeMuX_1_4_st
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY DeMuX_1_4_TB IS
END DeMuX_1_4_TB;
 
ARCHITECTURE behavior OF DeMuX_1_4_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT DeMuX_1_4_st
    PORT(
         a : IN  std_logic;
         s : IN  std_logic_vector(1 downto 0);
         z : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic := '0';
   signal s : std_logic_vector(1 downto 0) := (others => '0');

 	--Outputs
   signal z : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DeMuX_1_4_st PORT MAP (
          a => a,
          s => s,
          z => z
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

--      wait for <clock>_period*10;

      -- insert stimulus here 
		a <= '1';
		s(1) <= '0'; s(0) <= '0'; wait for 100 ns;
		s(1) <= '0'; s(0) <= '1'; wait for 100 ns;
		s(1) <= '1'; s(0) <= '0'; wait for 100 ns;
		s(1) <= '1'; s(0) <= '1'; wait for 100 ns;
      wait;
   end process;

END;
